module clockN(clk,q);
	input clk;
	output q;

	assign q = clk;

endmodule